* F:\CONTROL\COMPLMNT\CONVELV.SCH

* Schematics Version 6.1a - August 1994
* Thu Jan 28 13:52:21 1999


** Analysis setup **
.tran 10us 10ms
.OP 


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib nom.lib

.INC "CONVELV.net"
.INC "CONVELV.als"


.probe


.END
